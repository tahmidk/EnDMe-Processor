/**---------------------------------------------------------------------
 *	Module:		Top Level EnDMe Processor
 *	Class:		CSE 141L - SP18
 * Authors: 	Tahmid Khan
 *					Shengyuan Lin
 *----------------------------------------------------------------------
 *	[Description]
 *	This module puts the EnDMe processor together module by module based
 * on the high level block diagram
 *
 *	[Input]
 *		CLK - the clock (1-bit)
 *		reset_ctrl - the control wire that resets pc to 0 if high (1-bit)
 *
 *	[Output]
 *		None - check that data_mem has correct outputs
 ---------------------------------------------------------------------*/
 
 module top_level(
	input CLK,
	input reset_ctrl
 );
 
	// Initialize instruction fetch
	instr_fetch IF(
	
	);
	
	// Initialize instruction ROM
	instr_rom IROM(
	
	);
	
	// Initialize ALU
	alu ALU(
	
	);
	
	// Initialize accumulator
	accumulator ACC(
	
	);
	
	// Initialize control unit
	
	// Initialize register file
	
	// Initialize data memory
	
	// Initialize
 
 
 endmodule